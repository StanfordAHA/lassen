// Stub impl until coreir supports bfloat verilog generation
module mul (
  input [15:0] in0,
  input [15:0] in1,
  output [15:0] out
);
assign out = 0;

endmodule
